module Ejer2(
  input isZero,
  input isBEQ,
  input isBNE,
  input isJmp,
  input [31:0] currentPC,
  input [31:0] jmpTarget32,
  input [31:0] branchTargetAddr,
  output [31:0] nextPC
);

  // TODO: Compute nextPC value

endmodule
